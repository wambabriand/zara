
module PIXEL #parameter( N = 8 ) (

		input [N:0] I ,
		input [N:0] O ,
		output  clk
) ;






endmodule 
