

module MED #(parameter N = 7, M = 8)(
 input [N:0]  DI, 
 input BYP,  clk, DSI ,
 output logic [N:0] D
) ;



wire [N:0] w0,w1,w2,w3,w4,w5,w6,w7 ;
int i;


always @(clk)

  begin

	for(i=0;i<M;i++){
		
	}
	


  end

endmodule
